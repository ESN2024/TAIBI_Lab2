
module TAIBI_Lab2 (
	clk_clk,
	digit_1_external_connection_export,
	reset_reset_n,
	start_external_connection_export);	

	input		clk_clk;
	output	[3:0]	digit_1_external_connection_export;
	input		reset_reset_n;
	input		start_external_connection_export;
endmodule
